module filterGPU ();



endmodule 