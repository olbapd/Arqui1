module dkSideMem(input logic [9:0]horz,vert,
					 output logic [2:0] draw_dk);
					 
	logic [0:2]RAM [0:31] [0:63] ='{'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b010,3'b011,3'b011,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b001,3'b001,3'b010,3'b010,3'b010,3'b011,3'b001,3'b010,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b001,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b001,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b010,3'b001,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b001,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b001,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b001,3'b010,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b001,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b001,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b001,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b010,3'b001,3'b010,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b010,3'b010,3'b001,3'b001,3'b010,3'b001,3'b001,3'b010,3'b001,3'b010,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000},
'{3'b000,3'b010,3'b010,3'b010,3'b001,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b010,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000}};
		
		
		logic [2:0] temp;
		assign temp	= RAM[vert][horz];
		always_comb begin 
			if (temp === 3'bxxx) begin
				draw_dk = 3'b000;
			end
			else begin 
				draw_dk = temp;

			end
		end
endmodule