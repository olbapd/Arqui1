module pizzaMem(input logic [9:0]horz,vert,
					 output logic [1:0] draw_pizza);
	logic [0:1]RAM [0:31] [0:31] ='{'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b01,2'b01,2'b01,2'b01,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b01,2'b01,2'b10,2'b10,2'b10,2'b01,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b01,2'b10,2'b10,2'b10,2'b01,2'b01,2'b01,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b01,2'b10,2'b10,2'b01,2'b01,2'b11,2'b11,2'b11,2'b01,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b01,2'b10,2'b10,2'b01,2'b11,2'b11,2'b11,2'b01,2'b01,2'b01,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b01,2'b10,2'b10,2'b01,2'b11,2'b11,2'b11,2'b01,2'b10,2'b10,2'b01,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b01,2'b10,2'b10,2'b01,2'b11,2'b11,2'b11,2'b11,2'b01,2'b10,2'b10,2'b01,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b01,2'b10,2'b01,2'b11,2'b01,2'b01,2'b11,2'b11,2'b11,2'b01,2'b01,2'b11,2'b01,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b01,2'b10,2'b10,2'b01,2'b01,2'b10,2'b10,2'b01,2'b11,2'b11,2'b11,2'b11,2'b11,2'b01,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b01,2'b10,2'b01,2'b11,2'b01,2'b10,2'b10,2'b01,2'b11,2'b11,2'b11,2'b11,2'b11,2'b01,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b01,2'b10,2'b01,2'b11,2'b11,2'b01,2'b01,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b01,2'b01,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b01,2'b01,2'b01,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b01,2'b01,2'b11,2'b11,2'b01,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b01,2'b01,2'b01,2'b01,2'b01,2'b11,2'b01,2'b10,2'b10,2'b01,2'b11,2'b01,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b01,2'b01,2'b01,2'b01,2'b10,2'b01,2'b11,2'b01,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b01,2'b01,2'b01,2'b01,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00},
'{2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00}};
		
		
		//assign draw_pizza = RAM[vert][horz];
		logic [1:0] temp;
		assign temp	= RAM[vert][horz];
		always_comb begin 
			if (temp === 2'bxx) begin
				draw_pizza = 2'b00;
			end
			else begin 
				draw_pizza = RAM[vert][horz];

			end
		end

endmodule
