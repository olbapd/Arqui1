module instrcutionMem 
			#(parameter N=32)
			(  input logic [N-1:0] addr,
				output logic [N-1:0] instr)
		
		/*logic RAM[]
		
		
		always_comb begin 
			instr <= 
				
		end*/

endmodule