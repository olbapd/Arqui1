import utils::*;

module hazard_unit (
    input decode_execute_t dec_exe,
    input execute_memory exe_mem,
    input memory_writeback mem_wb,
    output hazard_unit_signals hazars_signals
);
    
endmodule


