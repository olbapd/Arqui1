module DecodeTB ();

	logic clk, RegWriteW,ImmSrcD;
    logic [31:0] Instr;
    logic [2:0][17:0] wd3;
    logic [3:0] wa3w;
    logic [2:0] RegSrc;
    logic [2:0][17:0] rd1, rd2;
    logic [2:0][17:0] ExtImm;

	initial begin

	end

endmodule