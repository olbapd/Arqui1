import utils::*;

