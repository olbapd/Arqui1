module imem (
    input logic [31:0] pc,
    output logic [31:0] Instr );

logic [31:0] RAM[64:0];

initial

$readmemh("C://",RAM);

assign Instr = RAM[pc[31:2]]; // word aligned